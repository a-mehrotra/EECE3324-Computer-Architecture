`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Aryan Mehrotra
// 
// Module Name: ID_EX_DFF
// Description: D Flip-Flop from instruction decode to execute stage
// Project Name: Final Project
//////////////////////////////////////////////////////////////////////////////////


module ID_EX_DFF(

    );
endmodule
