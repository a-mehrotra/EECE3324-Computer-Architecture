`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Aryan Mehrotra
// 
// Module Name: cpu5arm
// Description: Top file for ARM LEGV8 CPU
// Project Name: Final Project
//////////////////////////////////////////////////////////////////////////////////


module cpu5arm(ibus, clk, reset, iaddrbus, daddrbus, databus);
    input [31:0] ibus;
    input clk, reset;
    output [63:0] iaddrbus, daddrbus, databus;
    
    
endmodule
