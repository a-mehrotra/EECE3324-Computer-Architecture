`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Sam Bolduc and Aryan Mehrotra
// 
// Module Name: Controller
// Project Name: Assignment 4
//////////////////////////////////////////////////////////////////////////////////

module controller(ibus, clk, Cin, Imm, S, Aselect, Bselect, Dselect);
    input[31:0] ibus;
    input clk;
    output[2:0] S;
    output Imm, Cin;
    output[31:0] Aselect, Bselect, Dselect;
    
    
    
endmodule
